/*------------------------------------------------------------------------------
 * File          : D_MEMORY.sv
 * Project       : RTL
 * Author        : epwebq
 * Creation date : Oct 20, 2025
 * Description   :
 *------------------------------------------------------------------------------*/

module D_MEMORY #() ();

endmodule