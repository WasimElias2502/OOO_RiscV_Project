/*------------------------------------------------------------------------------
 * File          : PROCESSOR_ENUM.svh
 * Project       : RTL
 * Author        : epwebq
 * Creation date : Jun 20, 2025
 * Description   :
 *------------------------------------------------------------------------------*/


//****************** Instruction Fetch Unit Enum *************************//

typedef enum {sb , uj , jalr , pc_plus_4} next_pc_t;


//****************** Reservation Station Unit Enum *************************//