`timescale 1ns/1ns

interface RS_SCHEDULER_IF;


endinterface