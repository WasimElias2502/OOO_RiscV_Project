

interface RS_SCHEDULER_IF;


endinterface